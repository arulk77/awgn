/*
 ROM file necessary for the logarithmic function
 */
module rom_log();
  endmodule